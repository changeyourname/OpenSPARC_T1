// ========== Copyright Header Begin ==========================================
// 
// OpenSPARC T1 Processor File: ddr_ch_b.v
// Copyright (c) 2006 Sun Microsystems, Inc.  All Rights Reserved.
// DO NOT ALTER OR REMOVE COPYRIGHT NOTICES.
// 
// The above named program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public
// License version 2 as published by the Free Software Foundation.
// 
// The above named program is distributed in the hope that it will be 
// useful, but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
// General Public License for more details.
// 
// You should have received a copy of the GNU General Public
// License along with this work; if not, write to the Free Software
// Foundation, Inc., 51 Franklin St, Fifth Floor, Boston, MA 02110-1301, USA.
// 
// ========== Copyright Header End ============================================
module ddr_ch_b(afo ,serial_in ,afi ,serial_out ,pad_clk_si ,testmode_l
      ,test_mode ,bypass_enable_out ,ps_select_out ,rclk ,se ,pad_clk_so
      ,update_dr_in ,dram_io_data_out ,spare_ddr_pin ,spare_ddr_data ,
     dram_io_ptr_clk_inv ,bso ,bsi ,bypass_enable_in ,mode_ctrl_out ,
     update_dr_out ,shift_dr_out ,clock_dr_out ,hiz_n_out ,ps_select_in
      ,mode_ctrl_in ,shift_dr_in ,clock_dr_in ,hiz_n_in ,strobe , arst_l_out,
     io_dram_data_in ,io_dram_ecc_in ,dram_io_addr ,dram_io_clk_enable ,
     dram_io_cke ,dram_io_bank ,dram_io_ras_l ,dram_io_write_en_l ,
     dram_io_cas_l ,dram_io_cs_l ,dram_dq ,dram_addr ,dram_cb ,dram_dqs
      ,dram_cke ,dram_ba ,dram_ck_n ,dram_ck_p ,io_dram_data_valid ,
     dram_ras_l ,dram_we_l ,dram_cas_l ,dram_cs_l ,burst_length_four ,
     dram_io_pad_clk_inv ,dram_io_pad_enable ,dram_io_drive_enable ,
     rst_l ,lpf_code ,dram_io_channel_disabled ,dram_io_drive_data ,cbu
      ,vdd_h ,cbd, dram_arst_l );
output [143:0]	afi ;
output [143:0]	serial_out ;
output [255:0]	io_dram_data_in ;
output [31:0]	io_dram_ecc_in ;
input [143:0]	afo ;
input [143:0]	serial_in ;
input [287:0]	dram_io_data_out ;
input [9:0]	spare_ddr_data ;
input [4:0]	dram_io_ptr_clk_inv ;
input [14:0]	dram_io_addr ;
input [2:0]	dram_io_bank ;
input [3:0]	dram_io_cs_l ;
input [4:0]	lpf_code ;
input [8:1]	cbu ;
input [8:1]	cbd ;
inout [9:0]	spare_ddr_pin ;
inout [127:0]	dram_dq ;
inout [14:0]	dram_addr ;
inout [15:0]	dram_cb ;
inout [35:0]	dram_dqs ;
inout [2:0]	dram_ba ;
inout [3:0]	dram_ck_n ;
inout [3:0]	dram_ck_p ;
inout [3:0]	dram_cs_l ;
output		arst_l_out ;
output		bypass_enable_out ;
output		ps_select_out ;
output		pad_clk_so ;
output		bso ;
output		mode_ctrl_out ;
output		update_dr_out ;
output		shift_dr_out ;
output		clock_dr_out ;
output		hiz_n_out ;
output		io_dram_data_valid ;
input		pad_clk_si ;
input		testmode_l ;
input		test_mode ;
input		rclk ;
input		se ;
input		update_dr_in ;
input		bsi ;
input		bypass_enable_in ;
input		ps_select_in ;
input		mode_ctrl_in ;
input		shift_dr_in ;
input		clock_dr_in ;
input		hiz_n_in ;
input		strobe ;
input		dram_io_clk_enable ;
input		dram_io_cke ;
input		dram_io_ras_l ;
input		dram_io_write_en_l ;
input		dram_io_cas_l ;
input		burst_length_four ;
input		dram_io_pad_clk_inv ;
input		dram_io_pad_enable ;
input		dram_io_drive_enable ;
input		rst_l ;
input		dram_arst_l ;
input		dram_io_channel_disabled ;
input		dram_io_drive_data ;
input		vdd_h ;
inout		dram_cke ;
inout		dram_ras_l ;
inout		dram_we_l ;
inout		dram_cas_l ;
 
wire [8:1]	cbd_l ;
wire [7:0]	net0187 ;
wire [7:0]	net0182 ;
wire [7:0]	net0186 ;
wire [7:0]	net0412 ;
wire [7:0]	net0413 ;
wire [8:1]	cbu_l ;
wire [1:0]	pad_pos_cnt ;
wire [1:0]	pad_neg_cnt ;
wire		net0173 ;
wire		net0200 ;
wire		net0201 ;
wire		net0202 ;
wire		net0300 ;
wire		net0203 ;
wire		net0301 ;
wire		net0302 ;
wire		net0204 ;
wire		net0303 ;
wire		net0205 ;
wire		net0304 ;
wire		net0305 ;
wire		net0306 ;
wire		net0253 ;
wire		net0254 ;
wire		bso0_bsi1 ;
wire		pad_clk_so0_plogic_si1 ;
wire		se_out ;
wire		net0241 ;
wire		net0247 ;
wire		net0249 ;
wire		net0191 ;
wire		net0192 ;
wire		net0193 ;
wire		net0212 ;
wire		net0194 ;
wire		net0213 ;
wire		net0195 ;
wire		net0196 ;
wire		net0197 ;
wire		net0198 ;
wire		net0316 ;
wire		net0199 ;
wire		pvt_so_top_si ;
wire		plogic_clk_so1_pad_si2 ;
 
 
bw_io_ddr_sig_top_b I0 (
     .vrefcode_i_l    ({net0182[0] ,net0182[1] ,net0182[2] ,net0182[3] ,
            net0182[4] ,net0182[5] ,net0182[6] ,net0182[7] } ),
     .vrefcode_i_r    ({net0182[0] ,net0182[1] ,net0182[2] ,net0182[3] ,
            net0182[4] ,net0182[5] ,net0182[6] ,net0182[7] } ),
     .afo             ({afo[71:0] } ),
     .serial_in       ({serial_in[71:0] } ),
     .serial_out      ({serial_out[71:0] } ),
     .afi             ({afi[71:0] } ),
     .cbu_o_l         ({cbu_l } ),
     .cbd_o_l         ({cbd_l } ),
     .lpf_code_i_r    ({lpf_code } ),
     .dram_io_ptr_clk_inv_i_r ({dram_io_ptr_clk_inv[1:0] } ),
     .pad_pos_cnt_i_r ({pad_pos_cnt } ),
     .pad_neg_cnt_i_r ({pad_neg_cnt } ),
     .cbu_i_r         ({net0412[0] ,net0412[1] ,net0412[2] ,net0412[3] ,
            net0412[4] ,net0412[5] ,net0412[6] ,net0412[7] } ),
     .cbd_i_r         ({net0413[0] ,net0413[1] ,net0413[2] ,net0413[3] ,
            net0413[4] ,net0413[5] ,net0413[6] ,net0413[7] } ),
     .cbu_o_r         ({net0186[0] ,net0186[1] ,net0186[2] ,net0186[3] ,
            net0186[4] ,net0186[5] ,net0186[6] ,net0186[7] } ),
     .cbd_o_r         ({net0187[0] ,net0187[1] ,net0187[2] ,net0187[3] ,
            net0187[4] ,net0187[5] ,net0187[6] ,net0187[7] } ),
     .spare_ddr_data  ({spare_ddr_data[9:8] } ),
     .lpf_code_i_l    ({lpf_code } ),
     .dram_io_ptr_clk_inv_i_l ({dram_io_ptr_clk_inv[1:0] } ),
     .cbd_i_l         ({net0413[0] ,net0413[1] ,net0413[2] ,net0413[3] ,
            net0413[4] ,net0413[5] ,net0413[6] ,net0413[7] } ),
     .spare_ddr_pin   ({spare_ddr_pin[9:8] } ),
     .dram_ck_n       ({dram_ck_n } ),
     .dram_ck_p       ({dram_ck_p } ),
     .dram_io_bank    ({dram_io_bank[2] } ),
     .dram_ba         ({dram_ba[2] } ),
     .pad_neg_cnt_i_l ({pad_neg_cnt } ),
     .cbu_i_l         ({net0412[0] ,net0412[1] ,net0412[2] ,net0412[3] ,
            net0412[4] ,net0412[5] ,net0412[6] ,net0412[7] } ),
     .dram_cb         ({dram_cb[7:0] } ),
     .pad_pos_cnt_i_l ({pad_pos_cnt } ),
     .se_o_l          (se_out ),
     .dram_io_drive_enable_o_l (net0316 ),
     .mode_ctrl_out   (net0306 ),
     .update_dr_out   (net0305 ),
     .shift_dr_out    (net0304 ),
     .clock_dr_out    (net0303 ),
     .hiz_n_out       (net0302 ),
     .bypass_enable_out (net0301 ),
     .ps_select_out   (net0300 ),
     .test_mode_i_r   (test_mode ),
     .strobe_i_r      (strobe ),
     .testmode_l_i_l  (testmode_l ),
     .burst_length_four_i_r (burst_length_four ),
     .dram_io_pad_enable_i_r (dram_io_pad_enable ),
     .dram_io_drive_enable_i_r (dram_io_drive_enable ),
     .rst_l_i_r       (rst_l ),
     .arst_l_i_r      (dram_arst_l ),
     .dram_io_channel_disabled_i_r (dram_io_channel_disabled ),
     .dram_io_drive_data_i_r (dram_io_drive_data ),
     .se_i_r          (se ),
     .mode_ctrl_i_r   (net0191 ),
     .shift_dr_i_r    (net0193 ),
     .clock_dr_i_r    (net0194 ),
     .hiz_n_i_r       (net0195 ),
     .update_dr_i_r   (net0192 ),
     .vdd_h           (vdd_h ),
     .strobe_i_l      (strobe ),
     .bypass_enable_i_l (net0203 ),
     .ps_select_i_r   (net0197 ),
     .ps_select_i_l   (net0204 ),
     .test_mode_i_l   (test_mode ),
     .testmode_l_i_r  (testmode_l ),
     .dram_io_pad_enable_i_l (dram_io_pad_enable ),
     .burst_length_four_i_l (burst_length_four ),
     .\dram_io_data_out[95] (dram_io_data_out[95] ),
     .\dram_io_data_out[94] (dram_io_data_out[94] ),
     .\dram_io_data_out[93] (dram_io_data_out[93] ),
     .\dram_io_data_out[92] (dram_io_data_out[92] ),
     .\dram_io_data_out[91] (dram_io_data_out[91] ),
     .\dram_io_data_out[90] (dram_io_data_out[90] ),
     .\dram_io_data_out[89] (dram_io_data_out[89] ),
     .\dram_io_data_out[88] (dram_io_data_out[88] ),
     .\dram_io_data_out[87] (dram_io_data_out[87] ),
     .\dram_io_data_out[86] (dram_io_data_out[86] ),
     .\dram_io_data_out[85] (dram_io_data_out[85] ),
     .\dram_io_data_out[84] (dram_io_data_out[84] ),
     .\dram_io_data_out[83] (dram_io_data_out[83] ),
     .\dram_io_data_out[82] (dram_io_data_out[82] ),
     .\dram_io_data_out[81] (dram_io_data_out[81] ),
     .\dram_io_data_out[80] (dram_io_data_out[80] ),
     .\dram_io_data_out[79] (dram_io_data_out[79] ),
     .\dram_io_data_out[78] (dram_io_data_out[78] ),
     .\dram_io_data_out[77] (dram_io_data_out[77] ),
     .\dram_io_data_out[76] (dram_io_data_out[76] ),
     .\dram_io_data_out[75] (dram_io_data_out[75] ),
     .\dram_io_data_out[74] (dram_io_data_out[74] ),
     .\dram_io_data_out[73] (dram_io_data_out[73] ),
     .\dram_io_data_out[72] (dram_io_data_out[72] ),
     .\dram_io_data_out[71] (dram_io_data_out[71] ),
     .\dram_io_data_out[70] (dram_io_data_out[70] ),
     .\dram_io_data_out[69] (dram_io_data_out[69] ),
     .\dram_io_data_out[68] (dram_io_data_out[68] ),
     .\dram_io_data_out[67] (dram_io_data_out[67] ),
     .\dram_io_data_out[66] (dram_io_data_out[66] ),
     .\dram_io_data_out[65] (dram_io_data_out[65] ),
     .\dram_io_data_out[64] (dram_io_data_out[64] ),
     .\dram_io_data_out[31] (dram_io_data_out[31] ),
     .\dram_io_data_out[30] (dram_io_data_out[30] ),
     .\dram_io_data_out[29] (dram_io_data_out[29] ),
     .\dram_io_data_out[28] (dram_io_data_out[28] ),
     .\dram_io_data_out[27] (dram_io_data_out[27] ),
     .\dram_io_data_out[26] (dram_io_data_out[26] ),
     .\dram_io_data_out[25] (dram_io_data_out[25] ),
     .\dram_io_data_out[24] (dram_io_data_out[24] ),
     .\dram_io_data_out[23] (dram_io_data_out[23] ),
     .\dram_io_data_out[22] (dram_io_data_out[22] ),
     .\dram_io_data_out[21] (dram_io_data_out[21] ),
     .\dram_io_data_out[20] (dram_io_data_out[20] ),
     .\dram_io_data_out[19] (dram_io_data_out[19] ),
     .\dram_io_data_out[18] (dram_io_data_out[18] ),
     .\dram_io_data_out[17] (dram_io_data_out[17] ),
     .\dram_io_data_out[16] (dram_io_data_out[16] ),
     .\dram_io_data_out[15] (dram_io_data_out[15] ),
     .\dram_io_data_out[14] (dram_io_data_out[14] ),
     .\dram_io_data_out[13] (dram_io_data_out[13] ),
     .\dram_io_data_out[12] (dram_io_data_out[12] ),
     .\dram_io_data_out[11] (dram_io_data_out[11] ),
     .\dram_io_data_out[10] (dram_io_data_out[10] ),
     .\dram_io_data_out[9] (dram_io_data_out[9] ),
     .\dram_io_data_out[8] (dram_io_data_out[8] ),
     .\dram_io_data_out[7] (dram_io_data_out[7] ),
     .\dram_io_data_out[6] (dram_io_data_out[6] ),
     .\dram_io_data_out[5] (dram_io_data_out[5] ),
     .\dram_io_data_out[4] (dram_io_data_out[4] ),
     .\dram_io_data_out[3] (dram_io_data_out[3] ),
     .\dram_io_data_out[2] (dram_io_data_out[2] ),
     .\dram_io_data_out[1] (dram_io_data_out[1] ),
     .\dram_io_data_out[0] (dram_io_data_out[0] ),
     .dram_io_channel_disabled_i_l (dram_io_channel_disabled ),
     .dram_io_drive_enable_i_l (dram_io_drive_enable ),
     .rclk            (rclk ),
     .\dram_io_data_out[175] (dram_io_data_out[175] ),
     .\dram_io_data_out[174] (dram_io_data_out[174] ),
     .\dram_io_data_out[173] (dram_io_data_out[173] ),
     .\dram_io_data_out[172] (dram_io_data_out[172] ),
     .\dram_io_data_out[171] (dram_io_data_out[171] ),
     .\dram_io_data_out[170] (dram_io_data_out[170] ),
     .\dram_io_data_out[169] (dram_io_data_out[169] ),
     .\dram_io_data_out[168] (dram_io_data_out[168] ),
     .\dram_io_data_out[167] (dram_io_data_out[167] ),
     .\dram_io_data_out[166] (dram_io_data_out[166] ),
     .\dram_io_data_out[165] (dram_io_data_out[165] ),
     .\dram_io_data_out[164] (dram_io_data_out[164] ),
     .\dram_io_data_out[163] (dram_io_data_out[163] ),
     .\dram_io_data_out[162] (dram_io_data_out[162] ),
     .\dram_io_data_out[161] (dram_io_data_out[161] ),
     .\dram_io_data_out[160] (dram_io_data_out[160] ),
     .\dram_io_data_out[159] (dram_io_data_out[159] ),
     .\dram_io_data_out[158] (dram_io_data_out[158] ),
     .\dram_io_data_out[157] (dram_io_data_out[157] ),
     .\dram_io_data_out[156] (dram_io_data_out[156] ),
     .\dram_io_data_out[155] (dram_io_data_out[155] ),
     .\dram_io_data_out[154] (dram_io_data_out[154] ),
     .\dram_io_data_out[153] (dram_io_data_out[153] ),
     .\dram_io_data_out[152] (dram_io_data_out[152] ),
     .\dram_io_data_out[151] (dram_io_data_out[151] ),
     .\dram_io_data_out[150] (dram_io_data_out[150] ),
     .\dram_io_data_out[149] (dram_io_data_out[149] ),
     .\dram_io_data_out[148] (dram_io_data_out[148] ),
     .\dram_io_data_out[147] (dram_io_data_out[147] ),
     .\dram_io_data_out[146] (dram_io_data_out[146] ),
     .\dram_io_data_out[145] (dram_io_data_out[145] ),
     .\dram_io_data_out[144] (dram_io_data_out[144] ),
     .\dram_io_data_out[279] (dram_io_data_out[279] ),
     .\dram_io_data_out[278] (dram_io_data_out[278] ),
     .\dram_io_data_out[277] (dram_io_data_out[277] ),
     .\dram_io_data_out[276] (dram_io_data_out[276] ),
     .\dram_io_data_out[275] (dram_io_data_out[275] ),
     .\dram_io_data_out[274] (dram_io_data_out[274] ),
     .\dram_io_data_out[273] (dram_io_data_out[273] ),
     .\dram_io_data_out[272] (dram_io_data_out[272] ),
     .\io_dram_data_in[223] (io_dram_data_in[223] ),
     .\io_dram_data_in[222] (io_dram_data_in[222] ),
     .\io_dram_data_in[221] (io_dram_data_in[221] ),
     .\io_dram_data_in[220] (io_dram_data_in[220] ),
     .\io_dram_data_in[219] (io_dram_data_in[219] ),
     .\io_dram_data_in[218] (io_dram_data_in[218] ),
     .\io_dram_data_in[217] (io_dram_data_in[217] ),
     .\io_dram_data_in[216] (io_dram_data_in[216] ),
     .\io_dram_data_in[215] (io_dram_data_in[215] ),
     .\io_dram_data_in[214] (io_dram_data_in[214] ),
     .\io_dram_data_in[213] (io_dram_data_in[213] ),
     .\io_dram_data_in[212] (io_dram_data_in[212] ),
     .\io_dram_data_in[211] (io_dram_data_in[211] ),
     .\io_dram_data_in[210] (io_dram_data_in[210] ),
     .\io_dram_data_in[209] (io_dram_data_in[209] ),
     .\io_dram_data_in[208] (io_dram_data_in[208] ),
     .\io_dram_data_in[207] (io_dram_data_in[207] ),
     .\io_dram_data_in[206] (io_dram_data_in[206] ),
     .\io_dram_data_in[205] (io_dram_data_in[205] ),
     .\io_dram_data_in[204] (io_dram_data_in[204] ),
     .\io_dram_data_in[203] (io_dram_data_in[203] ),
     .\io_dram_data_in[202] (io_dram_data_in[202] ),
     .\io_dram_data_in[201] (io_dram_data_in[201] ),
     .\io_dram_data_in[200] (io_dram_data_in[200] ),
     .\io_dram_data_in[199] (io_dram_data_in[199] ),
     .\io_dram_data_in[198] (io_dram_data_in[198] ),
     .\io_dram_data_in[197] (io_dram_data_in[197] ),
     .\io_dram_data_in[196] (io_dram_data_in[196] ),
     .\io_dram_data_in[195] (io_dram_data_in[195] ),
     .\io_dram_data_in[194] (io_dram_data_in[194] ),
     .\io_dram_data_in[193] (io_dram_data_in[193] ),
     .\io_dram_data_in[192] (io_dram_data_in[192] ),
     .\dram_io_data_out[135] (dram_io_data_out[135] ),
     .\dram_io_data_out[134] (dram_io_data_out[134] ),
     .\dram_io_data_out[133] (dram_io_data_out[133] ),
     .\dram_io_data_out[132] (dram_io_data_out[132] ),
     .\dram_io_data_out[131] (dram_io_data_out[131] ),
     .\dram_io_data_out[130] (dram_io_data_out[130] ),
     .\dram_io_data_out[129] (dram_io_data_out[129] ),
     .\dram_io_data_out[128] (dram_io_data_out[128] ),
     .\io_dram_ecc_in[23] (io_dram_ecc_in[23] ),
     .\io_dram_ecc_in[22] (io_dram_ecc_in[22] ),
     .\io_dram_ecc_in[21] (io_dram_ecc_in[21] ),
     .\io_dram_ecc_in[20] (io_dram_ecc_in[20] ),
     .\io_dram_ecc_in[19] (io_dram_ecc_in[19] ),
     .\io_dram_ecc_in[18] (io_dram_ecc_in[18] ),
     .\io_dram_ecc_in[17] (io_dram_ecc_in[17] ),
     .\io_dram_ecc_in[16] (io_dram_ecc_in[16] ),
     .\io_dram_ecc_in[7] (io_dram_ecc_in[7] ),
     .\io_dram_ecc_in[6] (io_dram_ecc_in[6] ),
     .\io_dram_ecc_in[5] (io_dram_ecc_in[5] ),
     .\io_dram_ecc_in[4] (io_dram_ecc_in[4] ),
     .\io_dram_ecc_in[3] (io_dram_ecc_in[3] ),
     .\io_dram_ecc_in[2] (io_dram_ecc_in[2] ),
     .\io_dram_ecc_in[1] (io_dram_ecc_in[1] ),
     .\io_dram_ecc_in[0] (io_dram_ecc_in[0] ),
     .\io_dram_data_in[159] (io_dram_data_in[159] ),
     .\io_dram_data_in[158] (io_dram_data_in[158] ),
     .\io_dram_data_in[157] (io_dram_data_in[157] ),
     .\io_dram_data_in[156] (io_dram_data_in[156] ),
     .\io_dram_data_in[155] (io_dram_data_in[155] ),
     .\io_dram_data_in[154] (io_dram_data_in[154] ),
     .\io_dram_data_in[153] (io_dram_data_in[153] ),
     .\io_dram_data_in[152] (io_dram_data_in[152] ),
     .\io_dram_data_in[151] (io_dram_data_in[151] ),
     .\io_dram_data_in[150] (io_dram_data_in[150] ),
     .\io_dram_data_in[149] (io_dram_data_in[149] ),
     .\io_dram_data_in[148] (io_dram_data_in[148] ),
     .\io_dram_data_in[147] (io_dram_data_in[147] ),
     .\io_dram_data_in[146] (io_dram_data_in[146] ),
     .\io_dram_data_in[145] (io_dram_data_in[145] ),
     .\io_dram_data_in[144] (io_dram_data_in[144] ),
     .\io_dram_data_in[143] (io_dram_data_in[143] ),
     .\io_dram_data_in[142] (io_dram_data_in[142] ),
     .\io_dram_data_in[141] (io_dram_data_in[141] ),
     .\io_dram_data_in[140] (io_dram_data_in[140] ),
     .\io_dram_data_in[139] (io_dram_data_in[139] ),
     .\io_dram_data_in[138] (io_dram_data_in[138] ),
     .\io_dram_data_in[137] (io_dram_data_in[137] ),
     .\io_dram_data_in[136] (io_dram_data_in[136] ),
     .\io_dram_data_in[135] (io_dram_data_in[135] ),
     .\io_dram_data_in[134] (io_dram_data_in[134] ),
     .\io_dram_data_in[133] (io_dram_data_in[133] ),
     .\io_dram_data_in[132] (io_dram_data_in[132] ),
     .\io_dram_data_in[131] (io_dram_data_in[131] ),
     .\io_dram_data_in[130] (io_dram_data_in[130] ),
     .\io_dram_data_in[129] (io_dram_data_in[129] ),
     .\io_dram_data_in[128] (io_dram_data_in[128] ),
     .\io_dram_data_in[31] (io_dram_data_in[31] ),
     .\io_dram_data_in[30] (io_dram_data_in[30] ),
     .\io_dram_data_in[29] (io_dram_data_in[29] ),
     .\io_dram_data_in[28] (io_dram_data_in[28] ),
     .\io_dram_data_in[27] (io_dram_data_in[27] ),
     .\io_dram_data_in[26] (io_dram_data_in[26] ),
     .\io_dram_data_in[25] (io_dram_data_in[25] ),
     .\io_dram_data_in[24] (io_dram_data_in[24] ),
     .\io_dram_data_in[23] (io_dram_data_in[23] ),
     .\io_dram_data_in[22] (io_dram_data_in[22] ),
     .\io_dram_data_in[21] (io_dram_data_in[21] ),
     .\io_dram_data_in[20] (io_dram_data_in[20] ),
     .\io_dram_data_in[19] (io_dram_data_in[19] ),
     .\io_dram_data_in[18] (io_dram_data_in[18] ),
     .\io_dram_data_in[17] (io_dram_data_in[17] ),
     .\io_dram_data_in[16] (io_dram_data_in[16] ),
     .\io_dram_data_in[15] (io_dram_data_in[15] ),
     .\io_dram_data_in[14] (io_dram_data_in[14] ),
     .\io_dram_data_in[13] (io_dram_data_in[13] ),
     .\io_dram_data_in[12] (io_dram_data_in[12] ),
     .\io_dram_data_in[11] (io_dram_data_in[11] ),
     .\io_dram_data_in[10] (io_dram_data_in[10] ),
     .\io_dram_data_in[9] (io_dram_data_in[9] ),
     .\io_dram_data_in[8] (io_dram_data_in[8] ),
     .\io_dram_data_in[7] (io_dram_data_in[7] ),
     .\io_dram_data_in[6] (io_dram_data_in[6] ),
     .\io_dram_data_in[5] (io_dram_data_in[5] ),
     .\io_dram_data_in[4] (io_dram_data_in[4] ),
     .\io_dram_data_in[3] (io_dram_data_in[3] ),
     .\io_dram_data_in[2] (io_dram_data_in[2] ),
     .\io_dram_data_in[1] (io_dram_data_in[1] ),
     .\io_dram_data_in[0] (io_dram_data_in[0] ),
     .pad_clk_so      (pad_clk_so0_plogic_si1 ),
     .pad_clk_si      (pvt_so_top_si ),
     .\dram_addr[9]   (dram_addr[9] ),
     .\dram_addr[8]   (dram_addr[8] ),
     .\dram_addr[7]   (dram_addr[7] ),
     .\dram_addr[6]   (dram_addr[6] ),
     .\dram_addr[5]   (dram_addr[5] ),
     .\dram_addr[4]   (dram_addr[4] ),
     .\dram_addr[3]   (dram_addr[3] ),
     .\dram_addr[2]   (dram_addr[2] ),
     .\dram_addr[1]   (dram_addr[1] ),
     .\dram_addr[0]   (dram_addr[0] ),
     .\dram_io_addr[9] (dram_io_addr[9] ),
     .\dram_io_addr[8] (dram_io_addr[8] ),
     .\dram_io_addr[7] (dram_io_addr[7] ),
     .\dram_io_addr[6] (dram_io_addr[6] ),
     .\dram_io_addr[5] (dram_io_addr[5] ),
     .\dram_io_addr[4] (dram_io_addr[4] ),
     .\dram_io_addr[3] (dram_io_addr[3] ),
     .\dram_io_addr[2] (dram_io_addr[2] ),
     .\dram_io_addr[1] (dram_io_addr[1] ),
     .\dram_io_addr[0] (dram_io_addr[0] ),
     .\dram_dqs[12]   (dram_dqs[12] ),
     .\dram_dqs[11]   (dram_dqs[11] ),
     .\dram_dqs[10]   (dram_dqs[10] ),
     .\dram_dqs[9]    (dram_dqs[9] ),
     .\dram_dqs[8]    (dram_dqs[8] ),
     .bso             (bso0_bsi1 ),
     .bsi             (bsi ),
     .dram_io_clk_enable (dram_io_clk_enable ),
     .\dram_addr[14]  (dram_addr[14] ),
     .\dram_addr[13]  (dram_addr[13] ),
     .\dram_addr[12]  (dram_addr[12] ),
     .\dram_addr[11]  (dram_addr[11] ),
     .dram_cke        (dram_cke ),
     .dram_io_cke     (dram_io_cke ),
     .\dram_io_addr[14] (dram_io_addr[14] ),
     .\dram_io_addr[13] (dram_io_addr[13] ),
     .\dram_io_addr[12] (dram_io_addr[12] ),
     .\dram_io_addr[11] (dram_io_addr[11] ),
     .\dram_dq[95]    (dram_dq[95] ),
     .\dram_dq[94]    (dram_dq[94] ),
     .\dram_dq[93]    (dram_dq[93] ),
     .\dram_dq[92]    (dram_dq[92] ),
     .\dram_dq[91]    (dram_dq[91] ),
     .\dram_dq[90]    (dram_dq[90] ),
     .\dram_dq[89]    (dram_dq[89] ),
     .\dram_dq[88]    (dram_dq[88] ),
     .\dram_dq[87]    (dram_dq[87] ),
     .\dram_dq[86]    (dram_dq[86] ),
     .\dram_dq[85]    (dram_dq[85] ),
     .\dram_dq[84]    (dram_dq[84] ),
     .\dram_dq[83]    (dram_dq[83] ),
     .\dram_dq[82]    (dram_dq[82] ),
     .\dram_dq[81]    (dram_dq[81] ),
     .\dram_dq[80]    (dram_dq[80] ),
     .\dram_dq[79]    (dram_dq[79] ),
     .\dram_dq[78]    (dram_dq[78] ),
     .\dram_dq[77]    (dram_dq[77] ),
     .\dram_dq[76]    (dram_dq[76] ),
     .\dram_dq[75]    (dram_dq[75] ),
     .\dram_dq[74]    (dram_dq[74] ),
     .\dram_dq[73]    (dram_dq[73] ),
     .\dram_dq[72]    (dram_dq[72] ),
     .\dram_dq[71]    (dram_dq[71] ),
     .\dram_dq[70]    (dram_dq[70] ),
     .\dram_dq[69]    (dram_dq[69] ),
     .\dram_dq[68]    (dram_dq[68] ),
     .\dram_dq[67]    (dram_dq[67] ),
     .\dram_dq[66]    (dram_dq[66] ),
     .\dram_dq[65]    (dram_dq[65] ),
     .\dram_dq[64]    (dram_dq[64] ),
     .\dram_dq[31]    (dram_dq[31] ),
     .\dram_dq[30]    (dram_dq[30] ),
     .\dram_dq[29]    (dram_dq[29] ),
     .\dram_dq[28]    (dram_dq[28] ),
     .\dram_dq[27]    (dram_dq[27] ),
     .\dram_dq[26]    (dram_dq[26] ),
     .\dram_dq[25]    (dram_dq[25] ),
     .\dram_dq[24]    (dram_dq[24] ),
     .\dram_dq[23]    (dram_dq[23] ),
     .\dram_dq[22]    (dram_dq[22] ),
     .\dram_dq[21]    (dram_dq[21] ),
     .\dram_dq[20]    (dram_dq[20] ),
     .\dram_dq[19]    (dram_dq[19] ),
     .\dram_dq[18]    (dram_dq[18] ),
     .\dram_dq[17]    (dram_dq[17] ),
     .\dram_dq[16]    (dram_dq[16] ),
     .\dram_dq[15]    (dram_dq[15] ),
     .\dram_dq[14]    (dram_dq[14] ),
     .\dram_dq[13]    (dram_dq[13] ),
     .\dram_dq[12]    (dram_dq[12] ),
     .\dram_dq[11]    (dram_dq[11] ),
     .\dram_dq[10]    (dram_dq[10] ),
     .\dram_dq[9]     (dram_dq[9] ),
     .\dram_dq[8]     (dram_dq[8] ),
     .\dram_dq[7]     (dram_dq[7] ),
     .\dram_dq[6]     (dram_dq[6] ),
     .\dram_dq[5]     (dram_dq[5] ),
     .\dram_dq[4]     (dram_dq[4] ),
     .\dram_dq[3]     (dram_dq[3] ),
     .\dram_dq[2]     (dram_dq[2] ),
     .\dram_dq[1]     (dram_dq[1] ),
     .\dram_dq[0]     (dram_dq[0] ),
     .\dram_dqs[3]    (dram_dqs[3] ),
     .\dram_dqs[2]    (dram_dqs[2] ),
     .\dram_dqs[1]    (dram_dqs[1] ),
     .\dram_dqs[0]    (dram_dqs[0] ),
     .\dram_dqs[21]   (dram_dqs[21] ),
     .\dram_dqs[20]   (dram_dqs[20] ),
     .\dram_dqs[19]   (dram_dqs[19] ),
     .\dram_dqs[18]   (dram_dqs[18] ),
     .\dram_dqs[17]   (dram_dqs[17] ),
     .\dram_dqs[30]   (dram_dqs[30] ),
     .\dram_dqs[29]   (dram_dqs[29] ),
     .\dram_dqs[28]   (dram_dqs[28] ),
     .\dram_dqs[27]   (dram_dqs[27] ),
     .rst_l_i_l       (rst_l ),
     .arst_l_i_l      (dram_arst_l ),
     .bypass_enable_i_r (net0196 ),
     .hiz_n_i_l       (net0202 ),
     .shift_dr_i_l    (net0200 ),
     .mode_ctrl_i_l   (net0198 ),
     .dram_io_drive_data_i_l (dram_io_drive_data ),
     .se_i_l          (se ),
     .update_dr_i_l   (net0199 ),
     .clock_dr_i_l    (net0201 ),
     .\io_dram_data_in[95] (io_dram_data_in[95] ),
     .\io_dram_data_in[94] (io_dram_data_in[94] ),
     .\io_dram_data_in[93] (io_dram_data_in[93] ),
     .\io_dram_data_in[92] (io_dram_data_in[92] ),
     .\io_dram_data_in[91] (io_dram_data_in[91] ),
     .\io_dram_data_in[90] (io_dram_data_in[90] ),
     .\io_dram_data_in[89] (io_dram_data_in[89] ),
     .\io_dram_data_in[88] (io_dram_data_in[88] ),
     .\io_dram_data_in[87] (io_dram_data_in[87] ),
     .\io_dram_data_in[86] (io_dram_data_in[86] ),
     .\io_dram_data_in[85] (io_dram_data_in[85] ),
     .\io_dram_data_in[84] (io_dram_data_in[84] ),
     .\io_dram_data_in[83] (io_dram_data_in[83] ),
     .\io_dram_data_in[82] (io_dram_data_in[82] ),
     .\io_dram_data_in[81] (io_dram_data_in[81] ),
     .\io_dram_data_in[80] (io_dram_data_in[80] ),
     .\io_dram_data_in[79] (io_dram_data_in[79] ),
     .\io_dram_data_in[78] (io_dram_data_in[78] ),
     .\io_dram_data_in[77] (io_dram_data_in[77] ),
     .\io_dram_data_in[76] (io_dram_data_in[76] ),
     .\io_dram_data_in[75] (io_dram_data_in[75] ),
     .\io_dram_data_in[74] (io_dram_data_in[74] ),
     .\io_dram_data_in[73] (io_dram_data_in[73] ),
     .\io_dram_data_in[72] (io_dram_data_in[72] ),
     .\io_dram_data_in[71] (io_dram_data_in[71] ),
     .\io_dram_data_in[70] (io_dram_data_in[70] ),
     .\io_dram_data_in[69] (io_dram_data_in[69] ),
     .\io_dram_data_in[68] (io_dram_data_in[68] ),
     .\io_dram_data_in[67] (io_dram_data_in[67] ),
     .\io_dram_data_in[66] (io_dram_data_in[66] ),
     .\io_dram_data_in[65] (io_dram_data_in[65] ),
     .\io_dram_data_in[64] (io_dram_data_in[64] ),
     .\dram_io_data_out[239] (dram_io_data_out[239] ),
     .\dram_io_data_out[238] (dram_io_data_out[238] ),
     .\dram_io_data_out[237] (dram_io_data_out[237] ),
     .\dram_io_data_out[236] (dram_io_data_out[236] ),
     .\dram_io_data_out[235] (dram_io_data_out[235] ),
     .\dram_io_data_out[234] (dram_io_data_out[234] ),
     .\dram_io_data_out[233] (dram_io_data_out[233] ),
     .\dram_io_data_out[232] (dram_io_data_out[232] ),
     .\dram_io_data_out[231] (dram_io_data_out[231] ),
     .\dram_io_data_out[230] (dram_io_data_out[230] ),
     .\dram_io_data_out[229] (dram_io_data_out[229] ),
     .\dram_io_data_out[228] (dram_io_data_out[228] ),
     .\dram_io_data_out[227] (dram_io_data_out[227] ),
     .\dram_io_data_out[226] (dram_io_data_out[226] ),
     .\dram_io_data_out[225] (dram_io_data_out[225] ),
     .\dram_io_data_out[224] (dram_io_data_out[224] ),
     .\dram_io_data_out[223] (dram_io_data_out[223] ),
     .\dram_io_data_out[222] (dram_io_data_out[222] ),
     .\dram_io_data_out[221] (dram_io_data_out[221] ),
     .\dram_io_data_out[220] (dram_io_data_out[220] ),
     .\dram_io_data_out[219] (dram_io_data_out[219] ),
     .\dram_io_data_out[218] (dram_io_data_out[218] ),
     .\dram_io_data_out[217] (dram_io_data_out[217] ),
     .\dram_io_data_out[216] (dram_io_data_out[216] ),
     .\dram_io_data_out[215] (dram_io_data_out[215] ),
     .\dram_io_data_out[214] (dram_io_data_out[214] ),
     .\dram_io_data_out[213] (dram_io_data_out[213] ),
     .\dram_io_data_out[212] (dram_io_data_out[212] ),
     .\dram_io_data_out[211] (dram_io_data_out[211] ),
     .\dram_io_data_out[210] (dram_io_data_out[210] ),
     .\dram_io_data_out[209] (dram_io_data_out[209] ),
     .\dram_io_data_out[208] (dram_io_data_out[208] ) );
bw_io_ddr_sig_bot_b I1 (
     .vrefcode_i_l    ({net0182[0] ,net0182[1] ,net0182[2] ,net0182[3] ,
            net0182[4] ,net0182[5] ,net0182[6] ,net0182[7] } ),
     .vrefcode_i_r    ({net0182[0] ,net0182[1] ,net0182[2] ,net0182[3] ,
            net0182[4] ,net0182[5] ,net0182[6] ,net0182[7] } ),
     .serial_in       ({serial_in[143:72] } ),
     .afo             ({afo[143:72] } ),
     .serial_out      ({serial_out[143:72] } ),
     .afi             ({afi[143:72] } ),
     .spare_ddr_data  ({spare_ddr_data[7:0] } ),
     .spare_ddr_pin   ({spare_ddr_pin[7:0] } ),
     .cbu_i_r         ({net0186[0] ,net0186[1] ,net0186[2] ,net0186[3] ,
            net0186[4] ,net0186[5] ,net0186[6] ,net0186[7] } ),
     .cbd_i_r         ({net0187[0] ,net0187[1] ,net0187[2] ,net0187[3] ,
            net0187[4] ,net0187[5] ,net0187[6] ,net0187[7] } ),
     .dram_io_ptr_clk_inv_i_l ({dram_io_ptr_clk_inv[1:0] } ),
     .arst_l_out      (arst_l_out ),
     .lpf_code_i_l    ({lpf_code } ),
     .pad_pos_cnt_i_l ({pad_pos_cnt } ),
     .pad_neg_cnt_i_l ({pad_neg_cnt } ),
     .dram_cs_l       ({dram_cs_l } ),
     .cbu_i_l         ({cbu_l } ),
     .dram_cb         ({dram_cb[15:8] } ),
     .pad_neg_cnt_i_r ({pad_neg_cnt } ),
     .dram_io_bank    ({dram_io_bank[1:0] } ),
     .dram_addr       ({dram_addr[10] } ),
     .lpf_code_i_r    ({lpf_code } ),
     .cbd_i_l         ({cbd_l } ),
     .dram_io_ptr_clk_inv_i_r ({dram_io_ptr_clk_inv[1:0] } ),
     .dram_io_cs_l    ({dram_io_cs_l } ),
     .dram_ba         ({dram_ba[1:0] } ),
     .dram_io_addr    ({dram_io_addr[10] } ),
     .pad_pos_cnt_i_r ({pad_pos_cnt } ),
     .ps_select_i_r   (net0212 ),
     .test_mode_i_l   (test_mode ),
     .testmode_l_i_r  (testmode_l ),
     .test_mode_i_r   (test_mode ),
     .bypass_enable_i_l (net0213 ),
     .bypass_enable_i_r (net0213 ),
     .ps_select_i_l   (net0212 ),
     .update_dr_o_l   (net0199 ),
     .shift_dr_o_l    (net0200 ),
     .clock_dr_o_l    (net0201 ),
     .hiz_n_o_l       (net0202 ),
     .bypass_enable_o_l (net0203 ),
     .ps_select_o_r   (net0197 ),
     .mode_ctrl_o_r   (net0191 ),
     .update_dr_o_r   (net0192 ),
     .se_i_r          (se ),
     .mode_ctrl_i_r   (net0249 ),
     .clock_dr_i_r    (net0241 ),
     .mode_ctrl_o_l   (net0198 ),
     .hiz_n_i_r       (net0247 ),
     .update_dr_i_r   (net0254 ),
     .shift_dr_o_r    (net0193 ),
     .dram_io_drive_enable_i_r (dram_io_drive_enable ),
     .clock_dr_o_r    (net0194 ),
     .hiz_n_o_r       (net0195 ),
     .ps_select_o_l   (net0204 ),
     .rclk            (rclk ),
     .testmode_l_i_l  (testmode_l ),
     .burst_length_four_i_l (burst_length_four ),
     .dram_io_pad_enable_i_l (dram_io_pad_enable ),
     .dram_io_drive_enable_i_l (dram_io_drive_enable ),
     .rst_l_i_l       (rst_l ),
     .arst_l_i_l      (dram_arst_l ),
     .strobe_i_l      (strobe ),
     .dram_io_channel_disabled_i_l (dram_io_channel_disabled ),
     .dram_io_drive_data_i_l (dram_io_drive_data ),
     .dram_io_channel_disabled_i_r (dram_io_channel_disabled ),
     .dram_io_write_en_l (dram_io_write_en_l ),
     .\dram_io_data_out[63] (dram_io_data_out[63] ),
     .\dram_io_data_out[62] (dram_io_data_out[62] ),
     .\dram_io_data_out[61] (dram_io_data_out[61] ),
     .\dram_io_data_out[60] (dram_io_data_out[60] ),
     .\dram_io_data_out[59] (dram_io_data_out[59] ),
     .\dram_io_data_out[58] (dram_io_data_out[58] ),
     .\dram_io_data_out[57] (dram_io_data_out[57] ),
     .\dram_io_data_out[56] (dram_io_data_out[56] ),
     .\dram_io_data_out[55] (dram_io_data_out[55] ),
     .\dram_io_data_out[54] (dram_io_data_out[54] ),
     .\dram_io_data_out[53] (dram_io_data_out[53] ),
     .\dram_io_data_out[52] (dram_io_data_out[52] ),
     .\dram_io_data_out[51] (dram_io_data_out[51] ),
     .\dram_io_data_out[50] (dram_io_data_out[50] ),
     .\dram_io_data_out[49] (dram_io_data_out[49] ),
     .\dram_io_data_out[48] (dram_io_data_out[48] ),
     .\dram_io_data_out[47] (dram_io_data_out[47] ),
     .\dram_io_data_out[46] (dram_io_data_out[46] ),
     .\dram_io_data_out[45] (dram_io_data_out[45] ),
     .\dram_io_data_out[44] (dram_io_data_out[44] ),
     .\dram_io_data_out[43] (dram_io_data_out[43] ),
     .\dram_io_data_out[42] (dram_io_data_out[42] ),
     .\dram_io_data_out[41] (dram_io_data_out[41] ),
     .\dram_io_data_out[40] (dram_io_data_out[40] ),
     .\dram_io_data_out[39] (dram_io_data_out[39] ),
     .\dram_io_data_out[38] (dram_io_data_out[38] ),
     .\dram_io_data_out[37] (dram_io_data_out[37] ),
     .\dram_io_data_out[36] (dram_io_data_out[36] ),
     .\dram_io_data_out[35] (dram_io_data_out[35] ),
     .\dram_io_data_out[34] (dram_io_data_out[34] ),
     .\dram_io_data_out[33] (dram_io_data_out[33] ),
     .\dram_io_data_out[32] (dram_io_data_out[32] ),
     .\io_dram_data_in[255] (io_dram_data_in[255] ),
     .\io_dram_data_in[254] (io_dram_data_in[254] ),
     .\io_dram_data_in[253] (io_dram_data_in[253] ),
     .\io_dram_data_in[252] (io_dram_data_in[252] ),
     .\io_dram_data_in[251] (io_dram_data_in[251] ),
     .\io_dram_data_in[250] (io_dram_data_in[250] ),
     .\io_dram_data_in[249] (io_dram_data_in[249] ),
     .\io_dram_data_in[248] (io_dram_data_in[248] ),
     .\io_dram_data_in[247] (io_dram_data_in[247] ),
     .\io_dram_data_in[246] (io_dram_data_in[246] ),
     .\io_dram_data_in[245] (io_dram_data_in[245] ),
     .\io_dram_data_in[244] (io_dram_data_in[244] ),
     .\io_dram_data_in[243] (io_dram_data_in[243] ),
     .\io_dram_data_in[242] (io_dram_data_in[242] ),
     .\io_dram_data_in[241] (io_dram_data_in[241] ),
     .\io_dram_data_in[240] (io_dram_data_in[240] ),
     .\io_dram_data_in[239] (io_dram_data_in[239] ),
     .\io_dram_data_in[238] (io_dram_data_in[238] ),
     .\io_dram_data_in[237] (io_dram_data_in[237] ),
     .\io_dram_data_in[236] (io_dram_data_in[236] ),
     .\io_dram_data_in[235] (io_dram_data_in[235] ),
     .\io_dram_data_in[234] (io_dram_data_in[234] ),
     .\io_dram_data_in[233] (io_dram_data_in[233] ),
     .\io_dram_data_in[232] (io_dram_data_in[232] ),
     .\io_dram_data_in[231] (io_dram_data_in[231] ),
     .\io_dram_data_in[230] (io_dram_data_in[230] ),
     .\io_dram_data_in[229] (io_dram_data_in[229] ),
     .\io_dram_data_in[228] (io_dram_data_in[228] ),
     .\io_dram_data_in[227] (io_dram_data_in[227] ),
     .\io_dram_data_in[226] (io_dram_data_in[226] ),
     .\io_dram_data_in[225] (io_dram_data_in[225] ),
     .\io_dram_data_in[224] (io_dram_data_in[224] ),
     .dram_io_cas_l   (dram_io_cas_l ),
     .dram_we_l       (dram_we_l ),
     .dram_cas_l      (dram_cas_l ),
     .\dram_dq[127]   (dram_dq[127] ),
     .\dram_dq[126]   (dram_dq[126] ),
     .\dram_dq[125]   (dram_dq[125] ),
     .\dram_dq[124]   (dram_dq[124] ),
     .\dram_dq[123]   (dram_dq[123] ),
     .\dram_dq[122]   (dram_dq[122] ),
     .\dram_dq[121]   (dram_dq[121] ),
     .\dram_dq[120]   (dram_dq[120] ),
     .\dram_dq[119]   (dram_dq[119] ),
     .\dram_dq[118]   (dram_dq[118] ),
     .\dram_dq[117]   (dram_dq[117] ),
     .\dram_dq[116]   (dram_dq[116] ),
     .\dram_dq[115]   (dram_dq[115] ),
     .\dram_dq[114]   (dram_dq[114] ),
     .\dram_dq[113]   (dram_dq[113] ),
     .\dram_dq[112]   (dram_dq[112] ),
     .\dram_dq[111]   (dram_dq[111] ),
     .\dram_dq[110]   (dram_dq[110] ),
     .\dram_dq[109]   (dram_dq[109] ),
     .\dram_dq[108]   (dram_dq[108] ),
     .\dram_dq[107]   (dram_dq[107] ),
     .\dram_dq[106]   (dram_dq[106] ),
     .\dram_dq[105]   (dram_dq[105] ),
     .\dram_dq[104]   (dram_dq[104] ),
     .\dram_dq[103]   (dram_dq[103] ),
     .\dram_dq[102]   (dram_dq[102] ),
     .\dram_dq[101]   (dram_dq[101] ),
     .\dram_dq[100]   (dram_dq[100] ),
     .\dram_dq[99]    (dram_dq[99] ),
     .\dram_dq[98]    (dram_dq[98] ),
     .\dram_dq[97]    (dram_dq[97] ),
     .\dram_dq[96]    (dram_dq[96] ),
     .\dram_io_data_out[287] (dram_io_data_out[287] ),
     .\dram_io_data_out[286] (dram_io_data_out[286] ),
     .\dram_io_data_out[285] (dram_io_data_out[285] ),
     .\dram_io_data_out[284] (dram_io_data_out[284] ),
     .\dram_io_data_out[283] (dram_io_data_out[283] ),
     .\dram_io_data_out[282] (dram_io_data_out[282] ),
     .\dram_io_data_out[281] (dram_io_data_out[281] ),
     .\dram_io_data_out[280] (dram_io_data_out[280] ),
     .\dram_io_data_out[143] (dram_io_data_out[143] ),
     .\dram_io_data_out[142] (dram_io_data_out[142] ),
     .\dram_io_data_out[141] (dram_io_data_out[141] ),
     .\dram_io_data_out[140] (dram_io_data_out[140] ),
     .\dram_io_data_out[139] (dram_io_data_out[139] ),
     .\dram_io_data_out[138] (dram_io_data_out[138] ),
     .\dram_io_data_out[137] (dram_io_data_out[137] ),
     .\dram_io_data_out[136] (dram_io_data_out[136] ),
     .\io_dram_ecc_in[31] (io_dram_ecc_in[31] ),
     .\io_dram_ecc_in[30] (io_dram_ecc_in[30] ),
     .\io_dram_ecc_in[29] (io_dram_ecc_in[29] ),
     .\io_dram_ecc_in[28] (io_dram_ecc_in[28] ),
     .\io_dram_ecc_in[27] (io_dram_ecc_in[27] ),
     .\io_dram_ecc_in[26] (io_dram_ecc_in[26] ),
     .\io_dram_ecc_in[25] (io_dram_ecc_in[25] ),
     .\io_dram_ecc_in[24] (io_dram_ecc_in[24] ),
     .\io_dram_ecc_in[15] (io_dram_ecc_in[15] ),
     .\io_dram_ecc_in[14] (io_dram_ecc_in[14] ),
     .\io_dram_ecc_in[13] (io_dram_ecc_in[13] ),
     .\io_dram_ecc_in[12] (io_dram_ecc_in[12] ),
     .\io_dram_ecc_in[11] (io_dram_ecc_in[11] ),
     .\io_dram_ecc_in[10] (io_dram_ecc_in[10] ),
     .\io_dram_ecc_in[9] (io_dram_ecc_in[9] ),
     .\io_dram_ecc_in[8] (io_dram_ecc_in[8] ),
     .\dram_io_data_out[127] (dram_io_data_out[127] ),
     .\dram_io_data_out[126] (dram_io_data_out[126] ),
     .\dram_io_data_out[125] (dram_io_data_out[125] ),
     .\dram_io_data_out[124] (dram_io_data_out[124] ),
     .\dram_io_data_out[123] (dram_io_data_out[123] ),
     .\dram_io_data_out[122] (dram_io_data_out[122] ),
     .\dram_io_data_out[121] (dram_io_data_out[121] ),
     .\dram_io_data_out[120] (dram_io_data_out[120] ),
     .\dram_io_data_out[119] (dram_io_data_out[119] ),
     .\dram_io_data_out[118] (dram_io_data_out[118] ),
     .\dram_io_data_out[117] (dram_io_data_out[117] ),
     .\dram_io_data_out[116] (dram_io_data_out[116] ),
     .\dram_io_data_out[115] (dram_io_data_out[115] ),
     .\dram_io_data_out[114] (dram_io_data_out[114] ),
     .\dram_io_data_out[113] (dram_io_data_out[113] ),
     .\dram_io_data_out[112] (dram_io_data_out[112] ),
     .\dram_io_data_out[111] (dram_io_data_out[111] ),
     .\dram_io_data_out[110] (dram_io_data_out[110] ),
     .\dram_io_data_out[109] (dram_io_data_out[109] ),
     .\dram_io_data_out[108] (dram_io_data_out[108] ),
     .\dram_io_data_out[107] (dram_io_data_out[107] ),
     .\dram_io_data_out[106] (dram_io_data_out[106] ),
     .\dram_io_data_out[105] (dram_io_data_out[105] ),
     .\dram_io_data_out[104] (dram_io_data_out[104] ),
     .\dram_io_data_out[103] (dram_io_data_out[103] ),
     .\dram_io_data_out[102] (dram_io_data_out[102] ),
     .\dram_io_data_out[101] (dram_io_data_out[101] ),
     .\dram_io_data_out[100] (dram_io_data_out[100] ),
     .\dram_io_data_out[99] (dram_io_data_out[99] ),
     .\dram_io_data_out[98] (dram_io_data_out[98] ),
     .\dram_io_data_out[97] (dram_io_data_out[97] ),
     .\dram_io_data_out[96] (dram_io_data_out[96] ),
     .\io_dram_data_in[191] (io_dram_data_in[191] ),
     .\io_dram_data_in[190] (io_dram_data_in[190] ),
     .\io_dram_data_in[189] (io_dram_data_in[189] ),
     .\io_dram_data_in[188] (io_dram_data_in[188] ),
     .\io_dram_data_in[187] (io_dram_data_in[187] ),
     .\io_dram_data_in[186] (io_dram_data_in[186] ),
     .\io_dram_data_in[185] (io_dram_data_in[185] ),
     .\io_dram_data_in[184] (io_dram_data_in[184] ),
     .\io_dram_data_in[183] (io_dram_data_in[183] ),
     .\io_dram_data_in[182] (io_dram_data_in[182] ),
     .\io_dram_data_in[181] (io_dram_data_in[181] ),
     .\io_dram_data_in[180] (io_dram_data_in[180] ),
     .\io_dram_data_in[179] (io_dram_data_in[179] ),
     .\io_dram_data_in[178] (io_dram_data_in[178] ),
     .\io_dram_data_in[177] (io_dram_data_in[177] ),
     .\io_dram_data_in[176] (io_dram_data_in[176] ),
     .\io_dram_data_in[175] (io_dram_data_in[175] ),
     .\io_dram_data_in[174] (io_dram_data_in[174] ),
     .\io_dram_data_in[173] (io_dram_data_in[173] ),
     .\io_dram_data_in[172] (io_dram_data_in[172] ),
     .\io_dram_data_in[171] (io_dram_data_in[171] ),
     .\io_dram_data_in[170] (io_dram_data_in[170] ),
     .\io_dram_data_in[169] (io_dram_data_in[169] ),
     .\io_dram_data_in[168] (io_dram_data_in[168] ),
     .\io_dram_data_in[167] (io_dram_data_in[167] ),
     .\io_dram_data_in[166] (io_dram_data_in[166] ),
     .\io_dram_data_in[165] (io_dram_data_in[165] ),
     .\io_dram_data_in[164] (io_dram_data_in[164] ),
     .\io_dram_data_in[163] (io_dram_data_in[163] ),
     .\io_dram_data_in[162] (io_dram_data_in[162] ),
     .\io_dram_data_in[161] (io_dram_data_in[161] ),
     .\io_dram_data_in[160] (io_dram_data_in[160] ),
     .rst_l_i_r       (rst_l ),
     .arst_l_i_r      (dram_arst_l ),
     .\io_dram_data_in[127] (io_dram_data_in[127] ),
     .\io_dram_data_in[126] (io_dram_data_in[126] ),
     .\io_dram_data_in[125] (io_dram_data_in[125] ),
     .\io_dram_data_in[124] (io_dram_data_in[124] ),
     .\io_dram_data_in[123] (io_dram_data_in[123] ),
     .\io_dram_data_in[122] (io_dram_data_in[122] ),
     .\io_dram_data_in[121] (io_dram_data_in[121] ),
     .\io_dram_data_in[120] (io_dram_data_in[120] ),
     .\io_dram_data_in[119] (io_dram_data_in[119] ),
     .\io_dram_data_in[118] (io_dram_data_in[118] ),
     .\io_dram_data_in[117] (io_dram_data_in[117] ),
     .\io_dram_data_in[116] (io_dram_data_in[116] ),
     .\io_dram_data_in[115] (io_dram_data_in[115] ),
     .\io_dram_data_in[114] (io_dram_data_in[114] ),
     .\io_dram_data_in[113] (io_dram_data_in[113] ),
     .\io_dram_data_in[112] (io_dram_data_in[112] ),
     .\io_dram_data_in[111] (io_dram_data_in[111] ),
     .\io_dram_data_in[110] (io_dram_data_in[110] ),
     .\io_dram_data_in[109] (io_dram_data_in[109] ),
     .\io_dram_data_in[108] (io_dram_data_in[108] ),
     .\io_dram_data_in[107] (io_dram_data_in[107] ),
     .\io_dram_data_in[106] (io_dram_data_in[106] ),
     .\io_dram_data_in[105] (io_dram_data_in[105] ),
     .\io_dram_data_in[104] (io_dram_data_in[104] ),
     .\io_dram_data_in[103] (io_dram_data_in[103] ),
     .\io_dram_data_in[102] (io_dram_data_in[102] ),
     .\io_dram_data_in[101] (io_dram_data_in[101] ),
     .\io_dram_data_in[100] (io_dram_data_in[100] ),
     .\io_dram_data_in[99] (io_dram_data_in[99] ),
     .\io_dram_data_in[98] (io_dram_data_in[98] ),
     .\io_dram_data_in[97] (io_dram_data_in[97] ),
     .\io_dram_data_in[96] (io_dram_data_in[96] ),
     .pad_clk_si      (plogic_clk_so1_pad_si2 ),
     .dram_ras_l      (dram_ras_l ),
     .dram_io_pad_enable_i_r (dram_io_pad_enable ),
     .\dram_io_data_out[271] (dram_io_data_out[271] ),
     .\dram_io_data_out[270] (dram_io_data_out[270] ),
     .\dram_io_data_out[269] (dram_io_data_out[269] ),
     .\dram_io_data_out[268] (dram_io_data_out[268] ),
     .\dram_io_data_out[267] (dram_io_data_out[267] ),
     .\dram_io_data_out[266] (dram_io_data_out[266] ),
     .\dram_io_data_out[265] (dram_io_data_out[265] ),
     .\dram_io_data_out[264] (dram_io_data_out[264] ),
     .\dram_io_data_out[263] (dram_io_data_out[263] ),
     .\dram_io_data_out[262] (dram_io_data_out[262] ),
     .\dram_io_data_out[261] (dram_io_data_out[261] ),
     .\dram_io_data_out[260] (dram_io_data_out[260] ),
     .\dram_io_data_out[259] (dram_io_data_out[259] ),
     .\dram_io_data_out[258] (dram_io_data_out[258] ),
     .\dram_io_data_out[257] (dram_io_data_out[257] ),
     .\dram_io_data_out[256] (dram_io_data_out[256] ),
     .\dram_io_data_out[255] (dram_io_data_out[255] ),
     .\dram_io_data_out[254] (dram_io_data_out[254] ),
     .\dram_io_data_out[253] (dram_io_data_out[253] ),
     .\dram_io_data_out[252] (dram_io_data_out[252] ),
     .\dram_io_data_out[251] (dram_io_data_out[251] ),
     .\dram_io_data_out[250] (dram_io_data_out[250] ),
     .\dram_io_data_out[249] (dram_io_data_out[249] ),
     .\dram_io_data_out[248] (dram_io_data_out[248] ),
     .\dram_io_data_out[247] (dram_io_data_out[247] ),
     .\dram_io_data_out[246] (dram_io_data_out[246] ),
     .\dram_io_data_out[245] (dram_io_data_out[245] ),
     .\dram_io_data_out[244] (dram_io_data_out[244] ),
     .\dram_io_data_out[243] (dram_io_data_out[243] ),
     .\dram_io_data_out[242] (dram_io_data_out[242] ),
     .\dram_io_data_out[241] (dram_io_data_out[241] ),
     .\dram_io_data_out[240] (dram_io_data_out[240] ),
     .mode_ctrl_i_l   (net0249 ),
     .\dram_dqs[7]    (dram_dqs[7] ),
     .\dram_dqs[6]    (dram_dqs[6] ),
     .\dram_dqs[5]    (dram_dqs[5] ),
     .\dram_dqs[4]    (dram_dqs[4] ),
     .bsi             (bso0_bsi1 ),
     .bso             (bso_pre_latch ),
     .burst_length_four_i_r (burst_length_four ),
     .strobe_i_r      (strobe ),
     .update_dr_i_l   (net0254 ),
     .hiz_n_i_l       (net0247 ),
     .clock_dr_i_l    (net0241 ),
     .shift_dr_i_l    (net0253 ),
     .se_i_l          (se ),
     .pad_clk_so      (pad_clk_so ),
     .dram_io_ras_l   (dram_io_ras_l ),
     .\dram_dq[63]    (dram_dq[63] ),
     .\dram_dq[62]    (dram_dq[62] ),
     .\dram_dq[61]    (dram_dq[61] ),
     .\dram_dq[60]    (dram_dq[60] ),
     .\dram_dq[59]    (dram_dq[59] ),
     .\dram_dq[58]    (dram_dq[58] ),
     .\dram_dq[57]    (dram_dq[57] ),
     .\dram_dq[56]    (dram_dq[56] ),
     .\dram_dq[55]    (dram_dq[55] ),
     .\dram_dq[54]    (dram_dq[54] ),
     .\dram_dq[53]    (dram_dq[53] ),
     .\dram_dq[52]    (dram_dq[52] ),
     .\dram_dq[51]    (dram_dq[51] ),
     .\dram_dq[50]    (dram_dq[50] ),
     .\dram_dq[49]    (dram_dq[49] ),
     .\dram_dq[48]    (dram_dq[48] ),
     .\dram_dq[47]    (dram_dq[47] ),
     .\dram_dq[46]    (dram_dq[46] ),
     .\dram_dq[45]    (dram_dq[45] ),
     .\dram_dq[44]    (dram_dq[44] ),
     .\dram_dq[43]    (dram_dq[43] ),
     .\dram_dq[42]    (dram_dq[42] ),
     .\dram_dq[41]    (dram_dq[41] ),
     .\dram_dq[40]    (dram_dq[40] ),
     .\dram_dq[39]    (dram_dq[39] ),
     .\dram_dq[38]    (dram_dq[38] ),
     .\dram_dq[37]    (dram_dq[37] ),
     .\dram_dq[36]    (dram_dq[36] ),
     .\dram_dq[35]    (dram_dq[35] ),
     .\dram_dq[34]    (dram_dq[34] ),
     .\dram_dq[33]    (dram_dq[33] ),
     .\dram_dq[32]    (dram_dq[32] ),
     .\dram_dqs[35]   (dram_dqs[35] ),
     .\dram_dqs[34]   (dram_dqs[34] ),
     .\dram_dqs[33]   (dram_dqs[33] ),
     .\dram_dqs[32]   (dram_dqs[32] ),
     .\dram_dqs[31]   (dram_dqs[31] ),
     .\dram_dqs[16]   (dram_dqs[16] ),
     .\dram_dqs[15]   (dram_dqs[15] ),
     .\dram_dqs[14]   (dram_dqs[14] ),
     .\dram_dqs[13]   (dram_dqs[13] ),
     .\dram_dqs[26]   (dram_dqs[26] ),
     .\dram_dqs[25]   (dram_dqs[25] ),
     .\dram_dqs[24]   (dram_dqs[24] ),
     .\dram_dqs[23]   (dram_dqs[23] ),
     .\dram_dqs[22]   (dram_dqs[22] ),
     .dram_io_drive_data_i_r (dram_io_drive_data ),
     .shift_dr_i_r    (net0253 ),
     .bypass_enable_o_r (net0196 ),
     .vdd_h           (vdd_h ),
     .\io_dram_data_in[63] (io_dram_data_in[63] ),
     .\io_dram_data_in[62] (io_dram_data_in[62] ),
     .\io_dram_data_in[61] (io_dram_data_in[61] ),
     .\io_dram_data_in[60] (io_dram_data_in[60] ),
     .\io_dram_data_in[59] (io_dram_data_in[59] ),
     .\io_dram_data_in[58] (io_dram_data_in[58] ),
     .\io_dram_data_in[57] (io_dram_data_in[57] ),
     .\io_dram_data_in[56] (io_dram_data_in[56] ),
     .\io_dram_data_in[55] (io_dram_data_in[55] ),
     .\io_dram_data_in[54] (io_dram_data_in[54] ),
     .\io_dram_data_in[53] (io_dram_data_in[53] ),
     .\io_dram_data_in[52] (io_dram_data_in[52] ),
     .\io_dram_data_in[51] (io_dram_data_in[51] ),
     .\io_dram_data_in[50] (io_dram_data_in[50] ),
     .\io_dram_data_in[49] (io_dram_data_in[49] ),
     .\io_dram_data_in[48] (io_dram_data_in[48] ),
     .\io_dram_data_in[47] (io_dram_data_in[47] ),
     .\io_dram_data_in[46] (io_dram_data_in[46] ),
     .\io_dram_data_in[45] (io_dram_data_in[45] ),
     .\io_dram_data_in[44] (io_dram_data_in[44] ),
     .\io_dram_data_in[43] (io_dram_data_in[43] ),
     .\io_dram_data_in[42] (io_dram_data_in[42] ),
     .\io_dram_data_in[41] (io_dram_data_in[41] ),
     .\io_dram_data_in[40] (io_dram_data_in[40] ),
     .\io_dram_data_in[39] (io_dram_data_in[39] ),
     .\io_dram_data_in[38] (io_dram_data_in[38] ),
     .\io_dram_data_in[37] (io_dram_data_in[37] ),
     .\io_dram_data_in[36] (io_dram_data_in[36] ),
     .\io_dram_data_in[35] (io_dram_data_in[35] ),
     .\io_dram_data_in[34] (io_dram_data_in[34] ),
     .\io_dram_data_in[33] (io_dram_data_in[33] ),
     .\io_dram_data_in[32] (io_dram_data_in[32] ),
     .\dram_io_data_out[207] (dram_io_data_out[207] ),
     .\dram_io_data_out[206] (dram_io_data_out[206] ),
     .\dram_io_data_out[205] (dram_io_data_out[205] ),
     .\dram_io_data_out[204] (dram_io_data_out[204] ),
     .\dram_io_data_out[203] (dram_io_data_out[203] ),
     .\dram_io_data_out[202] (dram_io_data_out[202] ),
     .\dram_io_data_out[201] (dram_io_data_out[201] ),
     .\dram_io_data_out[200] (dram_io_data_out[200] ),
     .\dram_io_data_out[199] (dram_io_data_out[199] ),
     .\dram_io_data_out[198] (dram_io_data_out[198] ),
     .\dram_io_data_out[197] (dram_io_data_out[197] ),
     .\dram_io_data_out[196] (dram_io_data_out[196] ),
     .\dram_io_data_out[195] (dram_io_data_out[195] ),
     .\dram_io_data_out[194] (dram_io_data_out[194] ),
     .\dram_io_data_out[193] (dram_io_data_out[193] ),
     .\dram_io_data_out[192] (dram_io_data_out[192] ),
     .\dram_io_data_out[191] (dram_io_data_out[191] ),
     .\dram_io_data_out[190] (dram_io_data_out[190] ),
     .\dram_io_data_out[189] (dram_io_data_out[189] ),
     .\dram_io_data_out[188] (dram_io_data_out[188] ),
     .\dram_io_data_out[187] (dram_io_data_out[187] ),
     .\dram_io_data_out[186] (dram_io_data_out[186] ),
     .\dram_io_data_out[185] (dram_io_data_out[185] ),
     .\dram_io_data_out[184] (dram_io_data_out[184] ),
     .\dram_io_data_out[183] (dram_io_data_out[183] ),
     .\dram_io_data_out[182] (dram_io_data_out[182] ),
     .\dram_io_data_out[181] (dram_io_data_out[181] ),
     .\dram_io_data_out[180] (dram_io_data_out[180] ),
     .\dram_io_data_out[179] (dram_io_data_out[179] ),
     .\dram_io_data_out[178] (dram_io_data_out[178] ),
     .\dram_io_data_out[177] (dram_io_data_out[177] ),
     .\dram_io_data_out[176] (dram_io_data_out[176] ) );
dram_pad_logic I9 (
     .pad_neg_cnt     ({pad_neg_cnt } ),
     .pad_pos_cnt     ({pad_pos_cnt } ),
     .testmode_l      (testmode_l ),
     .pad_logic_clk_se (se ),
     .pad_logic_clk_si (pad_clk_so0_plogic_si1 ),
     .dram_io_pad_clk_inv (dram_io_pad_clk_inv ),
     .dram_io_pad_enable (dram_io_pad_enable ),
     .burst_length_four (burst_length_four ),
     .clk             (net0173 ),
     .io_dram_data_valid (io_dram_data_valid ),
     .arst_l           (dram_arst_l ),
     .rst_l            (rst_l ),
     .pad_logic_clk_so (plogic_clk_so1_pad_si2 ) );
bw_u1_buf_15x I140 (
     .z               (net0249 ),
     .a               (mode_ctrl_in ) );
bw_u1_buf_15x I141 (
     .z               (net0254 ),
     .a               (update_dr_in ) );
bw_u1_buf_15x I142 (
     .z               (net0253 ),
     .a               (shift_dr_in ) );
bw_u1_buf_15x I143 (
     .z               (net0241 ),
     .a               (clock_dr_in ) );
bw_u1_buf_15x I144 (
     .z               (net0247 ),
     .a               (hiz_n_in ) );
bw_u1_buf_15x I145 (
     .z               (net0213 ),
     .a               (bypass_enable_in ) );
bw_u1_buf_15x I146 (
     .z               (net0212 ),
     .a               (ps_select_in ) );
bw_u1_buf_15x I155 (
     .z               (shift_dr_out ),
     .a               (net0304 ) );
bw_u1_buf_15x I156 (
     .z               (mode_ctrl_out ),
     .a               (net0306 ) );
bw_u1_buf_15x I157 (
     .z               (bypass_enable_out ),
     .a               (net0301 ) );
bw_u1_buf_15x I158 (
     .z               (clock_dr_out ),
     .a               (net0303 ) );
bw_u1_buf_15x I159 (
     .z               (update_dr_out ),
     .a               (net0305 ) );
bw_u1_buf_15x I160 (
     .z               (hiz_n_out ),
     .a               (net0302 ) );
bw_u1_buf_15x I161 (
     .z               (ps_select_out ),
     .a               (net0300 ) );
bw_u1_buf_5x I172 (
     .z               (net0205 ),
     .a               (net0316 ) );
bw_io_ddr_pvt_enable I176 (
     .cbd_in          ({cbd } ),
     .cbu_in          ({cbu } ),
     .cbu_out         ({net0412[0] ,net0412[1] ,net0412[2] ,net0412[3] ,
            net0412[4] ,net0412[5] ,net0412[6] ,net0412[7] } ),
     .cbd_out         ({net0413[0] ,net0413[1] ,net0413[2] ,net0413[3] ,
            net0413[4] ,net0413[5] ,net0413[6] ,net0413[7] } ),
     .si              (pad_clk_si ),
     .en              (net0205 ),
     .rclk            (rclk ),
     .se              (se_out ),
     .so              (pvt_so_top_si ) );
bw_io_ddr_vref_logic I177 (
     .vrefcode        ({net0182[0] ,net0182[1] ,net0182[2] ,net0182[3] ,
            net0182[4] ,net0182[5] ,net0182[6] ,net0182[7] } ),
     .a               (dram_io_ptr_clk_inv[2] ),
     .c               (dram_io_ptr_clk_inv[4] ),
     .b               (dram_io_ptr_clk_inv[3] ),
     .vdd18           (vdd_h ) );
bw_u1_ckbuf_6x I124 (
     .clk             (net0173 ),
     .rclk            (rclk ) );
bw_u1_scanl_2x lockup_latch(
                .so(bso),
                .sd(bso_pre_latch),
                .ck(clock_dr_in));
endmodule
